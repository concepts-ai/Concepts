#!/usr/bin/env cdl-plan

problem "simple-float-csp"
domain "__empty__"

#!pragma load_implementation("3-simple-float-csp2.py")

def f(x: float32) -> float32

generator inv_f(x: float32, y: float32):
  goal: f(x) == y
  in: y
  out: x

generator inv_plus(x: float32, y: float32, z: float32):
  goal: x + y == z
  in: z, x
  out: y

generator gen_float(x: float32):
  out: x

controller print(s: string, x: float32)

behavior __goal__():
  body:
    bind x: float32
    bind y: float32

    assert f(x) + f(y) == 7.0
    print("x", x)
    print("y", y)

