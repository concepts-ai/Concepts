problem "blocksworld-sussman"
domain "blocksworld-breakdown.cdl"

#!pragma planner_is_goal_serializable=False
#!pragma planner_is_goal_ordered=True
#!pragma planner_always_commit_skeleton=True

objects:
  A: block
  B: block
  C: block

init:
  on_table[A] = True
  on_table[B] = True
  on[C, A] = True
  foreach x: block:
    clear[x] = True
  clear[A] = False
  handempty[...] = True


behavior __goal__():
  body:
    # Option 1
    foreach x: block:
      achieve_once on_table(x)

    # Option 2
    # foreach x: block:
    #   if not on_table(x):
    #     achieve_once on_table(x)

    # Option 3
    # achieve_once on_table(A)
    # achieve_once on_table(B)
    # achieve_once on_table(C)

    achieve_once handempty()

    achieve on(B, C)
    achieve on(A, B)
